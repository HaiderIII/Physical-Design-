// Module 1
module mod1(input a, output b);
endmodule
// Module 2
module mod2(input c, output d);
endmodule
// Module 3
module mod3(input e, output f);
endmodule
