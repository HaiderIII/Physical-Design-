// Module 2
module mod2(input c, output d);
endmodule
