module top (
    input clk,
    input rst,
    input [7:0] data_in,
    output [7:0] data_out
);

    wire w1, w2, w3;
    wire [7:0] internal_bus;
    reg [7:0] reg1, reg2;
    
    // Some logic here
    input signal1;
    input signal2;
    output result;
    
    wire temp1, temp2, temp3;
    
endmodule
