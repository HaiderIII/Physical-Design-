// Module 3
module mod3(input e, output f);
endmodule
