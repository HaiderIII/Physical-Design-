// Module 1
module mod1(input a, output b);
endmodule
